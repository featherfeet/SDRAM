// sdram_system_tb.v

// Generated using ACDS version 13.0sp1 232 at 2019.03.01.18:13:37

`timescale 1 ps / 1 ps
module sdram_system_tb (
	);

	wire         sdram_system_inst_clk_bfm_clk_clk;                            // sdram_system_inst_clk_bfm:clk -> [sdram_system_inst:clk_clk, sdram_system_inst_reset_bfm:clk]
	wire         sdram_system_inst_reset_bfm_reset_reset;                      // sdram_system_inst_reset_bfm:reset -> sdram_system_inst:reset_reset_n
	wire         sdram_system_inst_avalon_bridge_pins_acknowledge;             // sdram_system_inst:avalon_bridge_pins_acknowledge -> sdram_system_inst_avalon_bridge_pins_bfm:sig_acknowledge
	wire  [22:0] sdram_system_inst_avalon_bridge_pins_bfm_conduit_address;     // sdram_system_inst_avalon_bridge_pins_bfm:sig_address -> sdram_system_inst:avalon_bridge_pins_address
	wire  [15:0] sdram_system_inst_avalon_bridge_pins_read_data;               // sdram_system_inst:avalon_bridge_pins_read_data -> sdram_system_inst_avalon_bridge_pins_bfm:sig_read_data
	wire         sdram_system_inst_avalon_bridge_pins_bfm_conduit_write;       // sdram_system_inst_avalon_bridge_pins_bfm:sig_write -> sdram_system_inst:avalon_bridge_pins_write
	wire         sdram_system_inst_avalon_bridge_pins_bfm_conduit_read;        // sdram_system_inst_avalon_bridge_pins_bfm:sig_read -> sdram_system_inst:avalon_bridge_pins_read
	wire  [15:0] sdram_system_inst_avalon_bridge_pins_bfm_conduit_write_data;  // sdram_system_inst_avalon_bridge_pins_bfm:sig_write_data -> sdram_system_inst:avalon_bridge_pins_write_data
	wire   [1:0] sdram_system_inst_avalon_bridge_pins_bfm_conduit_byte_enable; // sdram_system_inst_avalon_bridge_pins_bfm:sig_byte_enable -> sdram_system_inst:avalon_bridge_pins_byte_enable
	wire         sdram_system_inst_sdram_controller_pins_cs_n;                 // sdram_system_inst:sdram_controller_pins_cs_n -> new_sdram_controller_0_my_partner:zs_cs_n
	wire   [1:0] sdram_system_inst_sdram_controller_pins_ba;                   // sdram_system_inst:sdram_controller_pins_ba -> new_sdram_controller_0_my_partner:zs_ba
	wire   [1:0] sdram_system_inst_sdram_controller_pins_dqm;                  // sdram_system_inst:sdram_controller_pins_dqm -> new_sdram_controller_0_my_partner:zs_dqm
	wire         sdram_system_inst_sdram_controller_pins_cke;                  // sdram_system_inst:sdram_controller_pins_cke -> new_sdram_controller_0_my_partner:zs_cke
	wire  [11:0] sdram_system_inst_sdram_controller_pins_addr;                 // sdram_system_inst:sdram_controller_pins_addr -> new_sdram_controller_0_my_partner:zs_addr
	wire         sdram_system_inst_sdram_controller_pins_we_n;                 // sdram_system_inst:sdram_controller_pins_we_n -> new_sdram_controller_0_my_partner:zs_we_n
	wire         sdram_system_inst_sdram_controller_pins_ras_n;                // sdram_system_inst:sdram_controller_pins_ras_n -> new_sdram_controller_0_my_partner:zs_ras_n
	wire         sdram_system_inst_sdram_controller_pins_cas_n;                // sdram_system_inst:sdram_controller_pins_cas_n -> new_sdram_controller_0_my_partner:zs_cas_n
	wire  [15:0] new_sdram_controller_0_my_partner_conduit_dq;                 // [] -> [new_sdram_controller_0_my_partner:zs_dq, sdram_system_inst:sdram_controller_pins_dq]
	wire         new_sdram_controller_0_my_partner_clk_bfm_clk_clk;            // new_sdram_controller_0_my_partner_clk_bfm:clk -> new_sdram_controller_0_my_partner:clk

	sdram_system sdram_system_inst (
		.clk_clk                        (sdram_system_inst_clk_bfm_clk_clk),                            //                   clk.clk
		.reset_reset_n                  (sdram_system_inst_reset_bfm_reset_reset),                      //                 reset.reset_n
		.sdram_controller_pins_addr     (sdram_system_inst_sdram_controller_pins_addr),                 // sdram_controller_pins.addr
		.sdram_controller_pins_ba       (sdram_system_inst_sdram_controller_pins_ba),                   //                      .ba
		.sdram_controller_pins_cas_n    (sdram_system_inst_sdram_controller_pins_cas_n),                //                      .cas_n
		.sdram_controller_pins_cke      (sdram_system_inst_sdram_controller_pins_cke),                  //                      .cke
		.sdram_controller_pins_cs_n     (sdram_system_inst_sdram_controller_pins_cs_n),                 //                      .cs_n
		.sdram_controller_pins_dq       (new_sdram_controller_0_my_partner_conduit_dq),                 //                      .dq
		.sdram_controller_pins_dqm      (sdram_system_inst_sdram_controller_pins_dqm),                  //                      .dqm
		.sdram_controller_pins_ras_n    (sdram_system_inst_sdram_controller_pins_ras_n),                //                      .ras_n
		.sdram_controller_pins_we_n     (sdram_system_inst_sdram_controller_pins_we_n),                 //                      .we_n
		.avalon_bridge_pins_address     (sdram_system_inst_avalon_bridge_pins_bfm_conduit_address),     //    avalon_bridge_pins.address
		.avalon_bridge_pins_byte_enable (sdram_system_inst_avalon_bridge_pins_bfm_conduit_byte_enable), //                      .byte_enable
		.avalon_bridge_pins_read        (sdram_system_inst_avalon_bridge_pins_bfm_conduit_read),        //                      .read
		.avalon_bridge_pins_write       (sdram_system_inst_avalon_bridge_pins_bfm_conduit_write),       //                      .write
		.avalon_bridge_pins_write_data  (sdram_system_inst_avalon_bridge_pins_bfm_conduit_write_data),  //                      .write_data
		.avalon_bridge_pins_acknowledge (sdram_system_inst_avalon_bridge_pins_acknowledge),             //                      .acknowledge
		.avalon_bridge_pins_read_data   (sdram_system_inst_avalon_bridge_pins_read_data)                //                      .read_data
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sdram_system_inst_clk_bfm (
		.clk (sdram_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sdram_system_inst_reset_bfm (
		.reset (sdram_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sdram_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm sdram_system_inst_avalon_bridge_pins_bfm (
		.sig_address     (sdram_system_inst_avalon_bridge_pins_bfm_conduit_address),     // conduit.address
		.sig_byte_enable (sdram_system_inst_avalon_bridge_pins_bfm_conduit_byte_enable), //        .byte_enable
		.sig_read        (sdram_system_inst_avalon_bridge_pins_bfm_conduit_read),        //        .read
		.sig_write       (sdram_system_inst_avalon_bridge_pins_bfm_conduit_write),       //        .write
		.sig_write_data  (sdram_system_inst_avalon_bridge_pins_bfm_conduit_write_data),  //        .write_data
		.sig_acknowledge (sdram_system_inst_avalon_bridge_pins_acknowledge),             //        .acknowledge
		.sig_read_data   (sdram_system_inst_avalon_bridge_pins_read_data)                //        .read_data
	);

	altera_sdram_partner_module new_sdram_controller_0_my_partner (
		.clk      (new_sdram_controller_0_my_partner_clk_bfm_clk_clk), //     clk.clk
		.zs_dq    (new_sdram_controller_0_my_partner_conduit_dq),      // conduit.dq
		.zs_addr  (sdram_system_inst_sdram_controller_pins_addr),      //        .addr
		.zs_ba    (sdram_system_inst_sdram_controller_pins_ba),        //        .ba
		.zs_cas_n (sdram_system_inst_sdram_controller_pins_cas_n),     //        .cas_n
		.zs_cke   (sdram_system_inst_sdram_controller_pins_cke),       //        .cke
		.zs_cs_n  (sdram_system_inst_sdram_controller_pins_cs_n),      //        .cs_n
		.zs_dqm   (sdram_system_inst_sdram_controller_pins_dqm),       //        .dqm
		.zs_ras_n (sdram_system_inst_sdram_controller_pins_ras_n),     //        .ras_n
		.zs_we_n  (sdram_system_inst_sdram_controller_pins_we_n)       //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) new_sdram_controller_0_my_partner_clk_bfm (
		.clk (new_sdram_controller_0_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
