// sdram_system.v

// Generated using ACDS version 13.0sp1 232 at 2019.03.01.18:13:47

`timescale 1 ps / 1 ps
module sdram_system (
		input  wire        clk_clk,                        //                   clk.clk
		input  wire        reset_reset_n,                  //                 reset.reset_n
		output wire [11:0] sdram_controller_pins_addr,     // sdram_controller_pins.addr
		output wire [1:0]  sdram_controller_pins_ba,       //                      .ba
		output wire        sdram_controller_pins_cas_n,    //                      .cas_n
		output wire        sdram_controller_pins_cke,      //                      .cke
		output wire        sdram_controller_pins_cs_n,     //                      .cs_n
		inout  wire [15:0] sdram_controller_pins_dq,       //                      .dq
		output wire [1:0]  sdram_controller_pins_dqm,      //                      .dqm
		output wire        sdram_controller_pins_ras_n,    //                      .ras_n
		output wire        sdram_controller_pins_we_n,     //                      .we_n
		input  wire [22:0] avalon_bridge_pins_address,     //    avalon_bridge_pins.address
		input  wire [1:0]  avalon_bridge_pins_byte_enable, //                      .byte_enable
		input  wire        avalon_bridge_pins_read,        //                      .read
		input  wire        avalon_bridge_pins_write,       //                      .write
		input  wire [15:0] avalon_bridge_pins_write_data,  //                      .write_data
		output wire        avalon_bridge_pins_acknowledge, //                      .acknowledge
		output wire [15:0] avalon_bridge_pins_read_data    //                      .read_data
	);

	wire         up_clocks_0_sdram_clk_clk;                                                 // up_clocks_0:SDRAM_CLK -> [bridge_0:clk, bridge_0_avalon_master_translator:clk, new_sdram_controller_0:clk, new_sdram_controller_0_s1_translator:clk, rst_controller_001:clk]
	wire         bridge_0_avalon_master_waitrequest;                                        // bridge_0_avalon_master_translator:av_waitrequest -> bridge_0:avalon_waitrequest
	wire  [22:0] bridge_0_avalon_master_address;                                            // bridge_0:avalon_address -> bridge_0_avalon_master_translator:av_address
	wire  [15:0] bridge_0_avalon_master_writedata;                                          // bridge_0:avalon_writedata -> bridge_0_avalon_master_translator:av_writedata
	wire         bridge_0_avalon_master_write;                                              // bridge_0:avalon_write -> bridge_0_avalon_master_translator:av_write
	wire         bridge_0_avalon_master_read;                                               // bridge_0:avalon_read -> bridge_0_avalon_master_translator:av_read
	wire  [15:0] bridge_0_avalon_master_readdata;                                           // bridge_0_avalon_master_translator:av_readdata -> bridge_0:avalon_readdata
	wire   [1:0] bridge_0_avalon_master_byteenable;                                         // bridge_0:avalon_byteenable -> bridge_0_avalon_master_translator:av_byteenable
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest;   // new_sdram_controller_0_s1_translator:uav_waitrequest -> bridge_0_avalon_master_translator:uav_waitrequest
	wire   [1:0] bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount;    // bridge_0_avalon_master_translator:uav_burstcount -> new_sdram_controller_0_s1_translator:uav_burstcount
	wire  [15:0] bridge_0_avalon_master_translator_avalon_universal_master_0_writedata;     // bridge_0_avalon_master_translator:uav_writedata -> new_sdram_controller_0_s1_translator:uav_writedata
	wire  [22:0] bridge_0_avalon_master_translator_avalon_universal_master_0_address;       // bridge_0_avalon_master_translator:uav_address -> new_sdram_controller_0_s1_translator:uav_address
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_lock;          // bridge_0_avalon_master_translator:uav_lock -> new_sdram_controller_0_s1_translator:uav_lock
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_write;         // bridge_0_avalon_master_translator:uav_write -> new_sdram_controller_0_s1_translator:uav_write
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_read;          // bridge_0_avalon_master_translator:uav_read -> new_sdram_controller_0_s1_translator:uav_read
	wire  [15:0] bridge_0_avalon_master_translator_avalon_universal_master_0_readdata;      // new_sdram_controller_0_s1_translator:uav_readdata -> bridge_0_avalon_master_translator:uav_readdata
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess;   // bridge_0_avalon_master_translator:uav_debugaccess -> new_sdram_controller_0_s1_translator:uav_debugaccess
	wire   [1:0] bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable;    // bridge_0_avalon_master_translator:uav_byteenable -> new_sdram_controller_0_s1_translator:uav_byteenable
	wire         bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid; // new_sdram_controller_0_s1_translator:uav_readdatavalid -> bridge_0_avalon_master_translator:uav_readdatavalid
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest;      // new_sdram_controller_0:za_waitrequest -> new_sdram_controller_0_s1_translator:av_waitrequest
	wire  [15:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata;        // new_sdram_controller_0_s1_translator:av_writedata -> new_sdram_controller_0:az_data
	wire  [21:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address;          // new_sdram_controller_0_s1_translator:av_address -> new_sdram_controller_0:az_addr
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect;       // new_sdram_controller_0_s1_translator:av_chipselect -> new_sdram_controller_0:az_cs
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write;            // new_sdram_controller_0_s1_translator:av_write -> new_sdram_controller_0:az_wr_n
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read;             // new_sdram_controller_0_s1_translator:av_read -> new_sdram_controller_0:az_rd_n
	wire  [15:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata;         // new_sdram_controller_0:za_data -> new_sdram_controller_0_s1_translator:av_readdata
	wire         new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid;    // new_sdram_controller_0:za_valid -> new_sdram_controller_0_s1_translator:av_readdatavalid
	wire   [1:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable;       // new_sdram_controller_0_s1_translator:av_byteenable -> new_sdram_controller_0:az_be_n
	wire         rst_controller_reset_out_reset;                                            // rst_controller:reset_out -> up_clocks_0:reset
	wire         rst_controller_001_reset_out_reset;                                        // rst_controller_001:reset_out -> [bridge_0:reset, bridge_0_avalon_master_translator:reset, new_sdram_controller_0:reset_n, new_sdram_controller_0_s1_translator:reset]

	sdram_system_up_clocks_0 up_clocks_0 (
		.CLOCK_50    (clk_clk),                        //       clk_in_primary.clk
		.reset       (rst_controller_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (),                               //              sys_clk.clk
		.sys_reset_n (),                               //        sys_clk_reset.reset_n
		.SDRAM_CLK   (up_clocks_0_sdram_clk_clk)       //            sdram_clk.clk
	);

	sdram_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (up_clocks_0_sdram_clk_clk),                                              //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                                    // reset.reset_n
		.az_addr        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_controller_pins_addr),                                             //  wire.export
		.zs_ba          (sdram_controller_pins_ba),                                               //      .export
		.zs_cas_n       (sdram_controller_pins_cas_n),                                            //      .export
		.zs_cke         (sdram_controller_pins_cke),                                              //      .export
		.zs_cs_n        (sdram_controller_pins_cs_n),                                             //      .export
		.zs_dq          (sdram_controller_pins_dq),                                               //      .export
		.zs_dqm         (sdram_controller_pins_dqm),                                              //      .export
		.zs_ras_n       (sdram_controller_pins_ras_n),                                            //      .export
		.zs_we_n        (sdram_controller_pins_we_n)                                              //      .export
	);

	sdram_system_bridge_0 bridge_0 (
		.clk                (up_clocks_0_sdram_clk_clk),          //        clock_reset.clk
		.reset              (rst_controller_001_reset_out_reset), //  clock_reset_reset.reset
		.avalon_readdata    (bridge_0_avalon_master_readdata),    //      avalon_master.readdata
		.avalon_waitrequest (bridge_0_avalon_master_waitrequest), //                   .waitrequest
		.avalon_byteenable  (bridge_0_avalon_master_byteenable),  //                   .byteenable
		.avalon_read        (bridge_0_avalon_master_read),        //                   .read
		.avalon_write       (bridge_0_avalon_master_write),       //                   .write
		.avalon_writedata   (bridge_0_avalon_master_writedata),   //                   .writedata
		.avalon_address     (bridge_0_avalon_master_address),     //                   .address
		.address            (avalon_bridge_pins_address),         // external_interface.export
		.byte_enable        (avalon_bridge_pins_byte_enable),     //                   .export
		.read               (avalon_bridge_pins_read),            //                   .export
		.write              (avalon_bridge_pins_write),           //                   .export
		.write_data         (avalon_bridge_pins_write_data),      //                   .export
		.acknowledge        (avalon_bridge_pins_acknowledge),     //                   .export
		.read_data          (avalon_bridge_pins_read_data)        //                   .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (23),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (23),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) bridge_0_avalon_master_translator (
		.clk                      (up_clocks_0_sdram_clk_clk),                                                 //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address              (bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (bridge_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (bridge_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (bridge_0_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (bridge_0_avalon_master_read),                                               //                          .read
		.av_readdata              (bridge_0_avalon_master_readdata),                                           //                          .readdata
		.av_write                 (bridge_0_avalon_master_write),                                              //                          .write
		.av_writedata             (bridge_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                          //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (23),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) new_sdram_controller_0_s1_translator (
		.clk                      (up_clocks_0_sdram_clk_clk),                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                    reset.reset
		.uav_address              (bridge_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (bridge_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read                 (bridge_0_avalon_master_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write                (bridge_0_avalon_master_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest          (bridge_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (bridge_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (bridge_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata             (bridge_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata            (bridge_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock                 (bridge_0_avalon_master_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess          (bridge_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.av_address               (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),          //      avalon_anti_slave_0.address
		.av_write                 (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),            //                         .write
		.av_read                  (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),             //                         .read
		.av_readdata              (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),         //                         .readdata
		.av_writedata             (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),        //                         .writedata
		.av_byteenable            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),       //                         .byteenable
		.av_readdatavalid         (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid),    //                         .readdatavalid
		.av_waitrequest           (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),      //                         .waitrequest
		.av_chipselect            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),       //                         .chipselect
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (up_clocks_0_sdram_clk_clk),          //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

endmodule
